typedef class eth_packet_chk_c ;
typedef class eth_packet_drv_c;
typedef class eth_packet_gen_c;
typedef class eth_packet_mon_c;
typedef class eth_packet_c;
typedef class packet_tb_env_c;
